int alu_passed_test_cases = 0; 
int alu_failed_test_cases = 0; 
static int  alu_golgen_output;