int top_passed_test_cases = 0; 
int top_failed_test_cases = 0; 
int golden_mux_out ; 