interface  top_intf;

    logic clk_top_intf;
    logic rst_top_intf; 
    logic sel_top_intf; 
    bit   [19:0] mux_out_top_intf; 
    
endinterface
