int reg_passed_test_cases = 0                ; 
int reg_failed_test_cases = 0                ; 
static reg [19:0] reg_golden_memory [15:0]   ; 
static int  reg_golgen_output                ;