int passed_test_cases;
int failed_test_cases;
bit [7:0] q_data; 
static int golden_P_Data; 
static int golden_Start; 
static int golden_parity; 
static int golden_end; 
static int golden_counter; 
int finish;