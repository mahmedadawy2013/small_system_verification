int reg2_passed_test_cases = 0; 
int reg2_failed_test_cases = 0; 
static reg [19:0] reg2_golden_memory [15:0]; 
static int  reg2_golgen_output;