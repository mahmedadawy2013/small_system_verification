
package pack1; 
    import uvm_pkg::*   ;
    `include "uvm_macros.svh"           
    `include "reg2_sequence_item.sv"
    `include "reg2_sequence.sv"
    `include "reg2_sequencer.sv"
    `include "reg2_driver.sv"   
    `include "reg2_monitor.sv"
    `include "reg2_agent_config.sv"
    `include "reg2_agent.sv"
    `include "reg2_scoreboard.sv"  
    `include "reg2_subscriber.sv" 
    `include "reg2_env_config.sv"
    `include "reg2_environment.sv"
    `include "reg2_test.sv"
endpackage 