
package pack1; 
    import uvm_pkg::*   ;
    `include "uvm_macros.svh"           
    `include "reg_sequence_item.sv"
    `include "reg_sequence.sv"
    `include "reg_sequencer.sv"
    `include "reg_driver.sv"   
    `include "reg_monitor.sv"
    `include "reg_agent_config.sv"
    `include "reg_agent.sv"
    `include "reg_scoreboard.sv"  
    `include "reg_subscriber.sv" 
    `include "reg_env_config.sv"
    `include "reg_environment.sv"
    `include "reg_test.sv"
    `include "reg_test_custoum.sv"
endpackage 