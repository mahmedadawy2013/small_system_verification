interface  top_intf;

    logic clk_top_intf;
    logic rst_top_intf; 
    logic sel_top_intf; 
    logic data_valid_top_intf;
    logic tx_out_top_intf;  
    logic busy_top_intf;    
    logic [19:0] mux_out_top_intf;
    
endinterface
